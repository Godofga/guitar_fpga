library verilog;
use verilog.vl_types.all;
entity teste0_vlg_vec_tst is
end teste0_vlg_vec_tst;
